io.phasetwo.keycloak.model.WebhookSpi
